// =============================================================================
// Module: gelu_unit
// Description: Combinational FP32 GeLU activation with a 256-entry LUT.
//              GeLU(x) = x * 0.5 * (1 + tanh(0.7978846*(x + 0.044715*x³)))
//              LUT covers x ∈ [-4.0, +3.96875], step 1/32 (addr = 128 + floor(x*32)).
//              x ≤ -4 → 0.0   |   x ≥ +4 → x (passthrough)   |   gelu_en=0 → bypass
//
// Generate gelu_lut.mem (run once before simulation/synthesis):
//   import struct, math
//   def fp32_hex(v): return '{:08x}'.format(struct.unpack('>I',struct.pack('>f',v))[0])
//   with open('gelu_lut.mem','w') as f:
//       for i in range(256):
//           x = max(-4.0, min(4.0, (i-128)/32.0))
//           g = x * 0.5 * (1 + math.tanh(0.7978846*(x + 0.044715*x**3)))
//           f.write(fp32_hex(g) + '\n')
// =============================================================================

module gelu_unit (
    input  logic [31:0] fp32_in,    // FP32 accumulator value
    input  logic        gelu_en,    // 1 = apply GeLU, 0 = bypass
    output logic [31:0] fp32_out    // FP32 GeLU(x) or x
);

    // =========================================================================
    // 256-entry FP32 LUT
    // Initialized from gelu_lut.mem (generated by the Python script above).
    // Each line is one 8-digit hex FP32 value, covering x = -4.0 to +3.96875.
    // =========================================================================
    logic [31:0] gelu_rom [0:255];
    initial $readmemh("gelu_lut.mem", gelu_rom);

    // =========================================================================
    // FP32 field extraction
    // =========================================================================
    logic        fp_sign;
    logic [7:0]  fp_exp;
    logic [22:0] fp_mant;

    assign fp_sign = fp32_in[31];
    assign fp_exp  = fp32_in[30:23];
    assign fp_mant = fp32_in[22:0];

    // abs_ge_4: |x| >= 4.0 (biased exp >= 129, covers NaN/Inf too)
    logic abs_ge_4;
    assign abs_ge_4 = (fp_exp >= 8'd129);

    // mag_idx = floor(|x| * 32) extracted from FP32 fields (no arithmetic needed).
    // Each biased exponent value shifts a different slice of the mantissa:
    //   exp=128 → [2,4): {1,   mant[22:17]}   exp=127 → [1,2): {01,  mant[22:18]}
    //   exp=126 → [.5,1):{001, mant[22:19]}   exp=125 → [.25,.5):{0001,mant[22:20]}
    //   exp=124 → [.125,.25):{00001,mant[22:21]}  exp=123 → [.0625,.125):{000001,mant[22]}
    //   exp<=122 or 0 → 0  (|x| < 0.0625 rounds to LUT entry at x=0)
    logic [6:0] mag_idx;

    always_comb begin
        case (fp_exp)
            8'd128: mag_idx = {1'b1,   fp_mant[22:17]};
            8'd127: mag_idx = {2'b01,  fp_mant[22:18]};
            8'd126: mag_idx = {3'b001, fp_mant[22:19]};
            8'd125: mag_idx = {4'b0001,fp_mant[22:20]};
            8'd124: mag_idx = {5'b00001,fp_mant[22:21]};
            8'd123: mag_idx = {6'b000001,fp_mant[22]};
            default: mag_idx = 7'd0;
        endcase
    end

    // LUT address: positive → 128 + mag_idx, negative → 128 - mag_idx
    logic [7:0] lut_addr;

    always_comb begin
        if (abs_ge_4)     lut_addr = 8'd0;
        else if (fp_sign) lut_addr = 8'd128 - {1'b0, mag_idx};
        else              lut_addr = 8'd128 + {1'b0, mag_idx};
    end

    always_comb begin
        if      (!gelu_en)              fp32_out = fp32_in;           // bypass
        else if (abs_ge_4 && fp_sign)   fp32_out = 32'h0000_0000;    // x <= -4 → 0
        else if (abs_ge_4 && !fp_sign)  fp32_out = fp32_in;          // x >= +4 → x
        else                            fp32_out = gelu_rom[lut_addr];
    end

endmodule
